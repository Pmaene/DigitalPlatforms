library ieee;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library work;
use work.std_logic_arithext.all;


-- datapath entity
entity my8051 is
port(
     RST                    : in  std_logic;
     CLK                    : in  std_logic
);
end my8051;


architecture RTL of my8051 is
begin

-- VHDL view of ipblock

end RTL;
